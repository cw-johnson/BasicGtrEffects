////////////////////////////////////////////////////////////////////////////	
//-------------------------------About------------------------------------// 
////////////////////////////////////////////////////////////////////////////
/*
Designer: Christopher Johnson
Graduate Project, DSP with FPGA's, Spring 2022
Professor Uwe Meyer-Baese
April 20, 2022





References and Credit
	The project used source code from Terasic's provided 'DE10_Standard_i2sound.v', and 'AUDIO_DAC.v'.
*/



//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module Basic_Gtr_Effects(

	//////////// CLOCK //////////
	input 		          		CLOCK2_50,
	input 		          		CLOCK3_50,
	input 		          		CLOCK4_50,
	input 		          		CLOCK_50,

	//////////// KEY //////////
	input 		     [3:0]		KEY,

	//////////// SW //////////
	input 		     [9:0]		SW,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// Seg7 //////////
	output		     [6:0]		HEX0,
	output		     [6:0]		HEX1,
	output		     [6:0]		HEX2,
	output		     [6:0]		HEX3,
	output		     [6:0]		HEX4,
	output		     [6:0]		HEX5,


	//////////// Audio //////////
	input		          		AUD_ADCDAT,
	input 		          		AUD_ADCLRCK,
	input 		          		AUD_BCLK,
	output	          		AUD_DACDAT,
	input 		          		AUD_DACLRCK,
	output		          		AUD_XCK,

	//////////// I2C for Audio and Video-In //////////
	output		          		FPGA_I2C_SCLK,
	inout 		          		FPGA_I2C_SDAT

);

////////////////////////////////////////////////////////////////////////////	
//----------------------I2C COdec Configuration---------------------------// 
////////////////////////////////////////////////////////////////////////////

//---------------------------------------------//
//-----I2C Message Transmit/Volume Control-----//
//---(From Terasic's de10_standard_i2sound.v)--//
//---------------------------------------------//
`define rom_size 7'd9  
parameter [8:0] DWIDTH = 8'd24;
parameter [8:0] AWIDTH = 8'd32;

reg  	[10:0]	COUNTER_500;
reg  	[15:0]	ROM[`rom_size-1:0];
reg  	[15:0]	DATA_A;
reg  	[5:0]	address;
wire CLOCK_500;
wire END;
wire KEY0_EDGE;
wire [23:0] DATA;
wire GO;
wire [3:0] level_vol;

assign CLOCK_500 = COUNTER_500[9]; //Clock/2^9=512
assign AUD_XCK 	= COUNTER_500[1]; //Clock/2^1=2
assign DATA = {8'h34, DATA_A};		//slave address + sub_address + register_data
assign GO = ((address <= `rom_size) && (END == 1)) ? COUNTER_500[10] : 1;


always @(posedge CLOCK_50) 
begin
	COUNTER_500=COUNTER_500+1;
end


always @(negedge KEY0_EDGE or posedge END) 
begin
	if (!KEY0_EDGE)
	begin
		address=0;
	end
	else if (address <= `rom_size)
	begin
		address=address+1;
	end
end

reg		[4:0]	vol;
wire	[6:0]	volume;

always @(negedge KEY0_EDGE or negedge KEY[1]) 
begin
	if(!KEY[1])
		vol = 5'd31;
	else if(vol == 5'd4)
		vol = 5'd31;
	else if(!KEY0_EDGE)
		vol = vol - 3;
end

//the volume level, level 0 to level 9,
//the higher the level, the greater the sound
assign level_vol = (vol - 4) / 3;
assign volume = vol + 96;

//--------------------------------------------------------//
//-------Parameterized WM8731 CODCEC Configuration ROM----//
//--------------------------------------------------------//
//Left Line In (0)
localparam LRINBOTH = 1'b0;
localparam LINMUTE = 1'b0;
localparam [4:0] LINVOL = 5'b10111;//0dB
//Right Line In (1)
localparam RLINBOTH = 1'b0;
localparam RINMUTE = 1'b1; //Mute
localparam [4:0] RINVOL = 5'b10111;//0dB
//Analogue Audio Path Control (4)
localparam [1:0] SIDEATT = 2'b00; //-6db
localparam SIDETONE = 1'b0; //Disable Sidetone
localparam DACSEL = 1'b1; //Select DAC
localparam BYPASS = 1'b0; //Disable Bypass
localparam INSEL = 1'b0; //Line in -> ADC
localparam MUTEMIC = 1'b1; //Mute Mic
localparam MICBOOST = 1'b0; //No Boost
//Digital Audio Path Control (5)
//Digital Audio Interface Format (7)
localparam BCLKINV = 1'b0; //Dont invert BCLK
localparam MS = 1'b1; //Master Mode
localparam LRSWAP = 1'b0; //Right DAC Data Right
localparam LRP = 1'b0; //Right channel DAC when DACLRC Low
localparam [1:0] IWL = 2'b10; //24 bits
localparam [1:0] FORMAT = 2'b10; //Left Justified I2S
//Sampling Control (8)
localparam CLKODIV2 = 1'b0; //Core Clock=CLOCKOUT
localparam CLKIDIV2 = 1'b0; //Core Clock=MCLK
localparam [3:0] SR = 4'b0111;
localparam BOSR = 1'b0; //256fs
localparam USBNORMAL = 1'b0; //Normal Mode

always @(posedge END) 
begin
	ROM[0] = {7'd0,LRINBOTH,LINMUTE,2'b00,LINVOL}; //Left Line In (0)
	ROM[1] = {7'd1,RLINBOTH,RINMUTE,2'b00,RINVOL}; //Right Line In (1)
	ROM[2] = {7'd2,2'b0,volume[6:0]};	//left channel headphone output volume
	ROM[3] = {7'd3,2'b0,volume[6:0]};	//right channel headphone output volume	
	ROM[4] = {7'd4,1'b0,SIDEATT,SIDETONE,DACSEL,BYPASS,INSEL,MUTEMIC,MICBOOST};
	ROM[5] = {7'd6,1'b0,8'h00}; //power down
	ROM[6] = {7'd7,1'b0,BCLKINV,MS,LRSWAP,LRP,IWL,FORMAT}; //Digital Audio Interface Format (7)
	ROM[7] = {7'd8,1'b0,CLKODIV2,CLKIDIV2,SR,BOSR,USBNORMAL}; //Sampling Control (8)
	ROM[8] = {7'd9,1'b0,8'h01};	//Active
	DATA_A = ROM[address];
end

//KEY trigger
keytr			u3(
	.clock(CLOCK_500),
	.key0(KEY[0]),
	.rst_n(KEY[1]),
	
	.KEY0_EDGE(KEY0_EDGE)
	);
				 
//i2c controller
i2c				u2( 
	// Host Side
	.CLOCK(CLOCK_500),
	.RESET(1'b1),
	// I2C Side
	.I2C_SDAT(FPGA_I2C_SDAT),
	.I2C_DATA(DATA),
	.I2C_SCLK(FPGA_I2C_SCLK),
	// Control Signals
	.GO(GO),
	.END(END)
	);
					 
HEX				u4(
	.hex(level_vol),
	.hex_fps(HEX0)
	);

HEX				u5(
	.hex({1'b0,GAIN1}),
	.hex_fps(HEX5)
	);	

HEX				u6(
	.hex({2'b00,CLIP}),
	.hex_fps(HEX4)
	);
	
HEX				u7(
	.hex({1'b0,FC}),
	.hex_fps(HEX3)
	);	
	
HEX				u8(
	.hex({1'b0,GAIN2}),
	.hex_fps(HEX2)
	);	
				
//--------------------------------------------------//	
//-------------Module Instantiation-----------------// 
//--------------------------------------------------//

wire signed [DWIDTH-1:0] I2S_AUDIO_IN, I2S_AUDIO_OUT;
wire signed [AWIDTH-1:0] GAIN1_AUDIO_IN, GAIN1_AUDIO_OUT;
wire signed [AWIDTH-1:0] SAT_AUDIO_IN, SAT_AUDIO_OUT;
wire signed [AWIDTH-1:0] LP_AUDIO_IN, LP_AUDIO_OUT;
wire signed [AWIDTH-1:0] GAIN2_AUDIO_IN, GAIN2_AUDIO_OUT;

wire [2:0] GAIN1, FC;
wire [2:0] GAIN2; 
wire [1:0] CLIP;
//Control Interface
assign GAIN1 = SW[2:0];
assign GAIN2 = {1'b0,SW[4:3]};
assign FC = SW[7:5];
assign CLIP = SW[9:8];

//Pipeline
//assign GAIN1_AUDIO_IN = $signed(I2S_AUDIO_OUT); //Sign Extend
//assign SAT_AUDIO_IN = GAIN1_AUDIO_OUT;
//assign LP_AUDIO_IN = SAT_AUDIO_OUT;
//assign GAIN2_AUDIO_IN = LP_AUDIO_OUT;
//assign I2S_AUDIO_IN = GAIN2_AUDIO_OUT >>> 8; //Discard Bits

assign GAIN1_AUDIO_IN = {{(AWIDTH-DWIDTH){I2S_AUDIO_OUT[23]}},I2S_AUDIO_OUT};//{I2S_AUDIO_OUT,8'd0}; //Sign Extend
assign SAT_AUDIO_IN = GAIN1_AUDIO_OUT;
assign LP_AUDIO_IN = SAT_AUDIO_OUT;
assign GAIN2_AUDIO_IN = LP_AUDIO_OUT;
assign I2S_AUDIO_IN = GAIN2_AUDIO_OUT; //Discard Bits

I2S_Interface #(DWIDTH) int0(AUD_BCLK,AUD_DACLRCK,AUD_ADCLRCK,AUD_DACDAT,AUD_ADCDAT,I2S_AUDIO_IN,I2S_AUDIO_OUT);

Gain_Stage #(AWIDTH) gain0(AUD_DACLRCK,GAIN1_AUDIO_IN,GAIN1_AUDIO_OUT,GAIN1);

Saturation_Stage #(AWIDTH) sat0(AUD_DACLRCK, SAT_AUDIO_IN, SAT_AUDIO_OUT, CLIP, LEDR[8],LEDR[9]);

IIR_LP_Filter #(AWIDTH) filt0(AUD_DACLRCK, LP_AUDIO_IN, LP_AUDIO_OUT, FC);

Gain_Stage #(AWIDTH) gain1(AUD_DACLRCK,GAIN2_AUDIO_IN,GAIN2_AUDIO_OUT,GAIN2);
//--------------------------------------------------//	
//---------------------Debugging--------------------// 
//--------------------------------------------------//
assign HEX1 = 7'h40;
assign LEDR[0] = GO;
assign LEDR[1] = END;
assign LEDR[2] = AUD_BCLK;
assign LEDR[3] = AUD_ADCLRCK;
assign LEDR[4] = AUD_DACLRCK;
assign LEDR[5] = AUD_ADCDAT;
assign LEDR[6] = AUD_DACDAT;
assign LEDR[7] = KEY0_EDGE;

endmodule	
	
	
	
	

	
	
//////////////////////////////////////////////////////////////////////////////	
//----------------------DAC I2S Interface/FSM-------------------------------// 
//////////////////////////////////////////////////////////////////////////////
module I2S_Interface
	#(parameter W = 24)(
	input BCLK, DACLRCK, ADCLRCK,
	output DACDAT, 
	input ADCDAT,
	input signed [W-1:0] AUDIO_IN,
	output reg signed [W-1:0] AUDIO_OUT
	);
	
localparam [4:0] S_STOP = 5'd24;
localparam [4:0] S_STANDBY = 5'd25;	
reg DACDAT_R;
reg [4:0] DAC_S, N_DAC_S, ADC_S, N_ADC_S;
reg signed [W-1:0] AUDIO_IN_BUF, AUDIO_OUT_BUF;	


initial begin
	DAC_S <= S_STANDBY; N_DAC_S <= S_STANDBY;	
	ADC_S <= S_STANDBY; N_DAC_S <= S_STANDBY;	
end


//DAC Next State Logic
always_comb begin
	if (DAC_S < W-1) //GO Transmit
		N_DAC_S <= DAC_S + 1'b1;
	else if (DAC_S == W-1)
		N_DAC_S <= S_STOP;
	else if (DAC_S == S_STOP)
		if (DACLRCK == 1'b1)
			N_DAC_S <= S_STANDBY;
		else
			N_DAC_S <= S_STOP;
	else if (DAC_S == S_STANDBY)
		if (DACLRCK == 1'b0)
			N_DAC_S <= 5'd0;
		else
			N_DAC_S <= S_STANDBY;
	else 
		N_DAC_S <= S_STOP;
end

//FSM Register
always @ (negedge BCLK) begin
	DAC_S <= N_DAC_S;
end

//DAC Output Logic
always_comb begin
	if (DAC_S < W)
		DACDAT_R <= AUDIO_OUT_BUF[W-1-DAC_S];
	else
		DACDAT_R <= 1'b0;
end
assign DACDAT = DACDAT_R;


//DAC FIFO Buffer
always @ (posedge DACLRCK) begin
	if (DACLRCK) begin
		AUDIO_OUT_BUF <= AUDIO_IN;
	end
end

////------------------ADC--------------------///
////ADC Next State Logic
always_comb begin
	if (ADC_S < W-1) //Go Recieve!
		N_ADC_S <= ADC_S + 1'b1;
	else if (ADC_S == W-1)
		N_ADC_S <= S_STOP;
	else if (ADC_S == S_STOP)
		if (ADCLRCK == 1'b1)
			N_ADC_S <= S_STANDBY;
		else
			N_ADC_S <= S_STOP;
	else if (ADC_S == S_STANDBY)
		if (ADCLRCK == 1'b0)
			N_ADC_S <= 5'd0;
		else
			N_ADC_S <= S_STANDBY;
	else 
		N_ADC_S <= S_STOP;
end

////FSM Register
always @ (negedge BCLK) begin
	ADC_S <= N_ADC_S;
	if (ADC_S < W)
		AUDIO_IN_BUF[W-1-ADC_S] <= ADCDAT;
end

////DAC FIFO Buffer
always @ (posedge DACLRCK)
	if (DACLRCK)
		AUDIO_OUT <= AUDIO_IN_BUF;

endmodule


//////////////////////////////////////////////////////////////////////////////	
//----------------------IIR Low-Pass Filter---------------------------------// 
//////////////////////////////////////////////////////////////////////////////
module IIR_LP_Filter
	#(parameter W = 32)(
	input DACLRCK,
	input signed [W-1:0] LP_IN,
	output reg signed [W-1:0] LP_OUT,
	input [3:0] FC
	);
////Low Pass Filter
wire signed [15:0] alpha = {8'd0,FC,4'd0};
wire signed [15:0] oneminalpha; 
assign oneminalpha =  16'b0000_0001_0000_0000 - alpha;
reg signed [47:0] LAST_Y, Y_LONG, X_LONG;

assign X_LONG = LP_IN <<< 8;
assign LP_OUT = Y_LONG >>> 9;
always @ (posedge DACLRCK) begin
	if (DACLRCK) begin
		Y_LONG <= X_LONG*alpha + LAST_Y*oneminalpha;
	end
end

endmodule



//////////////////////////////////////////////////////////////////////////////	
//-------------------------------Gain Stage---------------------------------// 
//////////////////////////////////////////////////////////////////////////////
module Gain_Stage
	#(parameter W = 32)(
	input DACLRCK,
	input signed [W-1:0] AUDIO_IN,
	output reg signed [W-1:0] AUDIO_OUT,
	input [2:0] GAIN_CONTROL
	);
	reg signed [7:0] GAIN;
	reg signed [W-1:0] res;

always_comb begin
	if (GAIN_CONTROL == 3'b000)
		GAIN <= 8'd0;
	else if (GAIN_CONTROL == 3'b001)
		GAIN <= 8'd1;
	else if (GAIN_CONTROL == 3'b010)
		GAIN <= 8'd2;
	else if (GAIN_CONTROL == 3'b011)
		GAIN <= 8'd4;
	else if (GAIN_CONTROL == 3'b100)
		GAIN <= 8'd8;
	else if (GAIN_CONTROL == 3'b101)
		GAIN <= 8'd16;
	else if (GAIN_CONTROL == 3'b110)
		GAIN <= 8'd32;
	else if (GAIN_CONTROL == 3'b111)
		GAIN <= 8'd64;
	else 
		GAIN <= 8'd0;
end

always @ (posedge DACLRCK) begin
	if (DACLRCK) begin
		AUDIO_OUT <= $signed(AUDIO_IN * GAIN) >>> 1;
	end
end
	
endmodule


//////////////////////////////////////////////////////////////////////////////	
//-------------------------Saturation Stage---------------------------------// 
//////////////////////////////////////////////////////////////////////////////
module Saturation_Stage
	#(parameter W = 32)(
	input DACLRCK,
	input signed[W-1:0] AUDIO_IN,
	output reg signed [W-1:0] AUDIO_OUT,
	input [1:0] saturation,
	output reg sat_debug1, sat_debug2
	);

localparam signed [W-1:0] T1 = 32'sd524_288;
localparam signed [W-1:0] T2 = 32'sd1_048_576;
localparam signed [W-1:0] T3 = 32'sd2_097_152;
reg signed [W-1:0] SAT_OUT1, SAT_OUT2, SAT_OUT3;

always @ (posedge DACLRCK) begin
	if (DACLRCK) begin
		AUDIO_OUT <= SAT_OUT3; //*AUDIO_IN*AUDIO_IN;
	end
end

always_comb begin
	if(AUDIO_IN > T1)
		sat_debug1 = 1'b1;
	else if(AUDIO_IN < -T1)
		sat_debug1 = 1'b1;	
	else
		sat_debug1 = 1'b0;
end

always_comb begin
	if(SAT_OUT1 > T2)
		sat_debug2 = 1'b1;
	else if(SAT_OUT1 < -T2)
		sat_debug2 = 1'b1;	
	else
		sat_debug2 = 1'b0;
end

always_comb begin
	if (saturation[0] == 1'b1) begin
		if (AUDIO_IN > T1) begin
			SAT_OUT1 <= T1 + (AUDIO_IN-T1)>>>1; 
		end else if (AUDIO_IN < -T1) begin
			SAT_OUT1 <= -T1 + (AUDIO_IN+T1)>>>1; 
		end else begin
			SAT_OUT1 <= AUDIO_IN; 
		end
	end else begin
		SAT_OUT1 <= AUDIO_IN;
	end
end

always_comb begin
	if (saturation[1] == 1'b1) begin
		if (SAT_OUT1 > T2) begin
			SAT_OUT2 <= T2 + (SAT_OUT1-T2)>>>2;; 
		end else if (SAT_OUT1 < -T2) begin
			SAT_OUT2 <= -T2 + (SAT_OUT1+T2)>>>2; 
		end else begin
			SAT_OUT2 <= SAT_OUT1; 
		end
	end else begin
		SAT_OUT2 <= SAT_OUT1;
	end
end

always_comb begin
	if (saturation == 2'b11) begin
		if (SAT_OUT2 > T3) begin
			SAT_OUT3 <= T3;
		end else if (SAT_OUT2 < -T3) begin
			SAT_OUT3 <= -T3; 
		end else begin
			SAT_OUT3 <= SAT_OUT2; 
		end
	end else begin
		SAT_OUT3 <= SAT_OUT2;
	end
end


endmodule





		

//////////////////////////////////////////////////////////////////////	
//--------------------------Sine Wave LUT ROM-----------------------// 
//////////////////////////////////////////////////////////////////////
module Sin_Gen(
	input DACLRCK,
	output signed [23:0] Sin_Gen_Out
	);
	
reg [7:0] SIN_Cont;
reg signed [15:0] Sin_Out;
assign Sin_Gen_Out = {Sin_Out,8'd0};

//Counter FSM
always @ (posedge DACLRCK) begin
	if (SIN_Cont < 47)
		SIN_Cont <= SIN_Cont + 1'b1;
	else 
		SIN_Cont <= 8'd0;
end

always@(SIN_Cont) begin
    case(SIN_Cont)
    0  :  Sin_Out       <=      0       ;
    1  :  Sin_Out       <=      4276    ;
    2  :  Sin_Out       <=      8480    ;
    3  :  Sin_Out       <=      12539   ;
    4  :  Sin_Out       <=      16383   ;
    5  :  Sin_Out       <=      19947   ;
    6  :  Sin_Out       <=      23169   ;
    7  :  Sin_Out       <=      25995   ;
    8  :  Sin_Out       <=      28377   ;
    9  :  Sin_Out       <=      30272   ;
    10  :  Sin_Out      <=      31650   ;
    11  :  Sin_Out      <=      32486   ;
    12  :  Sin_Out      <=      32767   ;
    13  :  Sin_Out      <=      32486   ;
    14  :  Sin_Out      <=      31650   ;
    15  :  Sin_Out      <=      30272   ;
    16  :  Sin_Out      <=      28377   ;
    17  :  Sin_Out      <=      25995   ;
    18  :  Sin_Out      <=      23169   ;
    19  :  Sin_Out      <=      19947   ;
    20  :  Sin_Out      <=      16383   ;
    21  :  Sin_Out      <=      12539   ;
    22  :  Sin_Out      <=      8480    ;
    23  :  Sin_Out      <=      4276    ;
    24  :  Sin_Out      <=      0       ;
    25  :  Sin_Out      <=      61259   ;
    26  :  Sin_Out      <=      57056   ;
    27  :  Sin_Out      <=      52997   ;
    28  :  Sin_Out      <=      49153   ;
    29  :  Sin_Out      <=      45589   ;
    30  :  Sin_Out      <=      42366   ;
    31  :  Sin_Out      <=      39540   ;
    32  :  Sin_Out      <=      37159   ;
    33  :  Sin_Out      <=      35263   ;
    34  :  Sin_Out      <=      33885   ;
    35  :  Sin_Out      <=      33049   ;
    36  :  Sin_Out      <=      32768   ;
    37  :  Sin_Out      <=      33049   ;
    38  :  Sin_Out      <=      33885   ;
    39  :  Sin_Out      <=      35263   ;
    40  :  Sin_Out      <=      37159   ;
    41  :  Sin_Out      <=      39540   ;
    42  :  Sin_Out      <=      42366   ;
    43  :  Sin_Out      <=      45589   ;
    44  :  Sin_Out      <=      49152   ;
    45  :  Sin_Out      <=      52997   ;
    46  :  Sin_Out      <=      57056   ;
    47  :  Sin_Out      <=      61259   ;
	default	:
		   Sin_Out		<=		0		;
	endcase
end
endmodule


